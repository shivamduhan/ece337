// $Id: $
// File name:   sensor_b.sv
// Created:     8/27/2019
// Author:      Shivam Duhan
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Behavorial style Sensor Error Detector Code
